module feedthru (
  input S,
  output Z
);

assign Z = S;

endmodule