.title <nem_ohmux_1b.sp>
.hdl nem_relay_1b.va

** Create relay and start at z=0 **
.subckt nem_ohmux_1b d s g b
    
.ends
** TODO! **
