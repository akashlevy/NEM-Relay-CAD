module feedthru (
  input I0,
  output Z
);

assign Z = I0;

endmodule