module feedthru (I0, Z);
  assign Z = I0;
endmodule